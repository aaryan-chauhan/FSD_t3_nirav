<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-9,15,113.4,-45.5</PageViewport>
<gate>
<ID>4</ID>
<type>AI_MUX_8x1</type>
<position>30,-17.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>10 </input>
<input>
<ID>IN_4</ID>11 </input>
<input>
<ID>IN_5</ID>12 </input>
<input>
<ID>IN_6</ID>13 </input>
<input>
<ID>IN_7</ID>14 </input>
<output>
<ID>OUT</ID>72 </output>
<input>
<ID>SEL_0</ID>3 </input>
<input>
<ID>SEL_1</ID>4 </input>
<input>
<ID>SEL_2</ID>2 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>25.5,-8.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>34.5,-8.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>30,-8</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>14,-28</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>14.5,-25</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>15,-22</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>16,-19</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>16,-16</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>15,-13.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>14.5,-10.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>13.5,-7.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AI_MUX_8x1</type>
<position>67.5,-20</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>50 </input>
<input>
<ID>IN_3</ID>51 </input>
<input>
<ID>IN_4</ID>50 </input>
<input>
<ID>IN_5</ID>51 </input>
<input>
<ID>IN_6</ID>51 </input>
<input>
<ID>IN_7</ID>50 </input>
<output>
<ID>OUT</ID>52 </output>
<input>
<ID>SEL_0</ID>48 </input>
<input>
<ID>SEL_1</ID>47 </input>
<input>
<ID>SEL_2</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>57</ID>
<type>AI_MUX_8x1</type>
<position>96,-20</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>53 </input>
<input>
<ID>IN_4</ID>55 </input>
<input>
<ID>IN_5</ID>53 </input>
<input>
<ID>IN_6</ID>53 </input>
<input>
<ID>IN_7</ID>53 </input>
<output>
<ID>OUT</ID>56 </output>
<input>
<ID>SEL_0</ID>49 </input>
<input>
<ID>SEL_1</ID>47 </input>
<input>
<ID>SEL_2</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>81,-3</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>81,-8</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>81,-11.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>77</ID>
<type>EE_VDD</type>
<position>51,-18.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>79</ID>
<type>FF_GND</type>
<position>51,-23.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>71.5,-20</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>EE_VDD</type>
<position>84,-18</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>85</ID>
<type>FF_GND</type>
<position>84,-21</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>100,-20</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_MUX_2x1</type>
<position>-57.5,-15.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>BA_DECODER_2x4</type>
<position>20,-48</position>
<input>
<ID>ENABLE</ID>61 </input>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT_0</ID>58 </output>
<output>
<ID>OUT_1</ID>57 </output>
<output>
<ID>OUT_2</ID>59 </output>
<output>
<ID>OUT_3</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>32.5,-48.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>60 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>11,-45</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>9.5,-48.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>11,-51</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>98</ID>
<type>AI_XOR2</type>
<position>85.5,-41</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AI_XOR2</type>
<position>85.5,-49</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AI_XOR2</type>
<position>85.5,-57</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>69,-37</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>69,-42</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>69,-50</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>69,-58</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>112</ID>
<type>GA_LED</type>
<position>89.5,-57</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>89.5,-41</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>89.5,-49</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>89.5,-34.5</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>GA_LED</type>
<position>34,-17.5</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-12,29,-11</points>
<connection>
<GID>4</GID>
<name>SEL_2</name></connection>
<intersection>-11 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25.5,-11,25.5,-10.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-11,29,-11</points>
<intersection>25.5 1</intersection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-12,31,-11</points>
<connection>
<GID>4</GID>
<name>SEL_0</name></connection>
<intersection>-11 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>34.5,-11,34.5,-10.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31,-11,34.5,-11</points>
<intersection>31 0</intersection>
<intersection>34.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-12,30,-10</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-12 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30,-12,30,-12</points>
<connection>
<GID>4</GID>
<name>SEL_1</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-28,22.5,-21</points>
<intersection>-28 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-21,27,-21</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-28,22.5,-28</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-25,21.5,-20</points>
<intersection>-25 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-20,27,-20</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-25,21.5,-25</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-22,20,-19</points>
<intersection>-22 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-19,27,-19</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-22,20,-22</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-18,27,-18</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>19 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>19,-19,19,-18</points>
<intersection>-19 8</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>18,-19,19,-19</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>19 4</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-17,27,-17</points>
<connection>
<GID>4</GID>
<name>IN_4</name></connection>
<intersection>19 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>19,-17,19,-16</points>
<intersection>-17 1</intersection>
<intersection>-16 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>18,-16,19,-16</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>19 5</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-16,20,-13.5</points>
<intersection>-16 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-16,27,-16</points>
<connection>
<GID>4</GID>
<name>IN_5</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-13.5,20,-13.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-15,21.5,-10.5</points>
<intersection>-15 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-15,27,-15</points>
<connection>
<GID>4</GID>
<name>IN_6</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-10.5,21.5,-10.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-14,22.5,-7.5</points>
<intersection>-14 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-14,27,-14</points>
<connection>
<GID>4</GID>
<name>IN_7</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-7.5,22.5,-7.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-14.5,67.5,-10</points>
<connection>
<GID>56</GID>
<name>SEL_1</name></connection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67.5,-10,96,-10</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>67.5 0</intersection>
<intersection>96 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>96,-14.5,96,-10</points>
<connection>
<GID>57</GID>
<name>SEL_1</name></connection>
<intersection>-10 2</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-14.5,95,-14</points>
<connection>
<GID>57</GID>
<name>SEL_2</name></connection>
<intersection>-14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>81,-14,81,-13.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-14,95,-14</points>
<intersection>68.5 4</intersection>
<intersection>81 1</intersection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>68.5,-14.5,68.5,-14</points>
<connection>
<GID>56</GID>
<name>SEL_0</name></connection>
<intersection>-14 2</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-14.5,97,-6</points>
<connection>
<GID>57</GID>
<name>SEL_0</name></connection>
<intersection>-6 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>81,-6,81,-5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-6,97,-6</points>
<intersection>66.5 4</intersection>
<intersection>81 1</intersection>
<intersection>97 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>66.5,-14.5,66.5,-6</points>
<connection>
<GID>56</GID>
<name>SEL_2</name></connection>
<intersection>-6 2</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-22.5,58,-16.5</points>
<intersection>-22.5 1</intersection>
<intersection>-21.5 6</intersection>
<intersection>-19.5 5</intersection>
<intersection>-18.5 2</intersection>
<intersection>-16.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-22.5,64.5,-22.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-18.5,58,-18.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>58,-16.5,64.5,-16.5</points>
<connection>
<GID>56</GID>
<name>IN_7</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>58,-19.5,64.5,-19.5</points>
<connection>
<GID>56</GID>
<name>IN_4</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>58,-21.5,64.5,-21.5</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-23.5,56,-17.5</points>
<intersection>-23.5 1</intersection>
<intersection>-20.5 7</intersection>
<intersection>-18.5 8</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-23.5,64.5,-23.5</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-17.5,64.5,-17.5</points>
<connection>
<GID>56</GID>
<name>IN_6</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>56,-20.5,64.5,-20.5</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>56,-18.5,64.5,-18.5</points>
<connection>
<GID>56</GID>
<name>IN_5</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-20,70.5,-20</points>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-20.5,89,-16.5</points>
<intersection>-20.5 2</intersection>
<intersection>-18.5 8</intersection>
<intersection>-18 1</intersection>
<intersection>-17.5 7</intersection>
<intersection>-16.5 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-18,89,-18</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-20.5,93,-20.5</points>
<connection>
<GID>57</GID>
<name>IN_3</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>89,-16.5,93,-16.5</points>
<connection>
<GID>57</GID>
<name>IN_7</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89,-17.5,93,-17.5</points>
<connection>
<GID>57</GID>
<name>IN_6</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89,-18.5,93,-18.5</points>
<connection>
<GID>57</GID>
<name>IN_5</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-23.5,87.5,-19.5</points>
<intersection>-23.5 1</intersection>
<intersection>-22.5 4</intersection>
<intersection>-21.5 5</intersection>
<intersection>-21 2</intersection>
<intersection>-19.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87.5,-23.5,93,-23.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-21,87.5,-21</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>87.5,-22.5,93,-22.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>87.5,-21.5,93,-21.5</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>87.5,-19.5,93,-19.5</points>
<connection>
<GID>57</GID>
<name>IN_4</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-20,99,-20</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<connection>
<GID>57</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-48.5,29.5,-48.5</points>
<connection>
<GID>90</GID>
<name>OUT_1</name></connection>
<connection>
<GID>92</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-49.5,29.5,-49.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-47.5,29.5,-47.5</points>
<connection>
<GID>90</GID>
<name>OUT_2</name></connection>
<connection>
<GID>92</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-46.5,29.5,-46.5</points>
<connection>
<GID>90</GID>
<name>OUT_3</name></connection>
<connection>
<GID>92</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-46.5,17,-45</points>
<connection>
<GID>90</GID>
<name>ENABLE</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-45,17,-45</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-51,14.5,-49.5</points>
<intersection>-51 2</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-49.5,17,-49.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-51,14.5,-51</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-48.5,17,-48.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-37,75,-37</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>75 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>75,-40,75,-34.5</points>
<intersection>-40 6</intersection>
<intersection>-37 1</intersection>
<intersection>-34.5 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>75,-40,82.5,-40</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>75 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>75,-34.5,88.5,-34.5</points>
<connection>
<GID>118</GID>
<name>N_in0</name></connection>
<intersection>75 4</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-42,82.5,-42</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>75 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>75,-48,75,-42</points>
<intersection>-48 5</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>75,-48,82.5,-48</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>75 4</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-50,82.5,-50</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>75 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75,-56,75,-50</points>
<intersection>-56 4</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>75,-56,82.5,-56</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>75 3</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-58,82.5,-58</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-49,88.5,-49</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<connection>
<GID>116</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-41,88.5,-41</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<connection>
<GID>114</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-57,88.5,-57</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>112</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-17.5,33,-17.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<connection>
<GID>122</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>